netcdf out {
dimensions:
	lat = 4 ;
	lon = 5 ;
variables:

	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:_CoordinateAxisType = "Lat" ;
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:_CoordinateAxisType = "Lon" ;

data:
     	lon=
       		10,15,20,25,30;
       	lat=	70,60,50,40;

group:  ROOT {
    variables:
         byte LAI(lat, lon) ;
         		LAI:CLASS = "DATA" ;
         		LAI:NB_BYTES = "Uint8" ;
         		LAI:_Unsigned = "true" ;
    data:
    	LAI=
    		20,20,20,30,30,
    		40,40,40,50,50,
    		60,60,60,70,70,
    		80,80,80,90,90;
    group: LEVEL1 {
        variables:
            byte V2(lat, lon) ;
                     		V2:CLASS = "DATA" ;
                     		V2:NB_BYTES = "Uint8" ;
                     		V2:_Unsigned = "true" ;
        data:
            	V2=
            		20,20,20,30,30,
            		40,40,40,50,50,
            		60,60,60,70,70,
            		80,80,80,90,90;
         }
    }
// global attributes:
		:_CoordSysBuilder = "ucar.nc2.dataset.conv.CF1Convention" ;
		:Conventions = "CF-1.5" ;


}
